vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|05 Sep 2011 17:02:23 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|05 Sep 2011 17:02:23 -0000
vti_filesize:IR|1419
vti_backlinkinfo:VX|
