vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|09 Feb 2014 13:25:45 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|09 Feb 2014 13:25:45 -0000
vti_filesize:IR|1039
vti_backlinkinfo:VX|
