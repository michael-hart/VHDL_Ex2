vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|06 Sep 2013 15:14:40 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|06 Sep 2013 15:14:40 -0000
vti_filesize:IR|4509
vti_backlinkinfo:VX|
